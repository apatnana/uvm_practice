//module tb;

//endmodule
